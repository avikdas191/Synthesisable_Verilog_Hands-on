module SevSeg(
	input  wire [3:0] HEX_2_disp,
	output wire [7:0] segments
);
	
	reg [7:0] tmp;
	
	always @(*)	begin
		case(HEX_2_disp)
			4'b0000: tmp = 8'b11000000;	// 0
			4'b0001: tmp = 8'b11111001;	// 1			
			4'b0010: tmp = 8'b10100100;	// 2
			4'b0011: tmp = 8'b10110000;	// 3
			4'b0100: tmp = 8'b10011001;	// 4			
			4'b0101: tmp = 8'b10010010;	// 5			
			4'b0110: tmp = 8'b10000010;	// 6
			4'b0111: tmp = 8'b11111000;	// 7			
			4'b1000: tmp = 8'b10000000;	// 8
			4'b1001: tmp = 8'b10010000;	// 9
			4'b1010: tmp = 8'b00001000;	// A			
			4'b1011: tmp = 8'b00000011;	// B
			4'b1100: tmp = 8'b01000110;	// C
			4'b1101: tmp = 8'b00100001;	// D			
			4'b1110: tmp = 8'b00000110;	// E
			4'b1111: tmp = 8'b00001110;	// F			
			default: tmp = 8'b11111111;	// blank - just in case
		endcase
	end

	assign segments = tmp;
	
endmodule
